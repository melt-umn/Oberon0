grammar edu:umn:cs:melt:Oberon0:core:concreteSyntax;

imports edu:umn:cs:melt:Oberon0:core:abstractSyntax;

imports silver:langutil only ast;

