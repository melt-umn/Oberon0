grammar edu:umn:cs:melt:Oberon0:constructs:dataStructures;

exports edu:umn:cs:melt:Oberon0:constructs:dataStructures:abstractSyntax;
exports edu:umn:cs:melt:Oberon0:constructs:dataStructures:concreteSyntax;

