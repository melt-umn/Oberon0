grammar edu:umn:cs:melt:Oberon0:constructs:procedures:concreteSyntax;

terminal Procedure_kwd 	'PROCEDURE' lexer classes {KEYWORD};


