grammar edu:umn:cs:melt:Oberon0:constructs:procedures:concreteSyntax;

imports silver:langutil:lsp as lsp;

terminal Procedure_kwd 	'PROCEDURE' lexer classes {KEYWORD};


