grammar edu:umn:cs:melt:Oberon0:components:L3;

exports edu:umn:cs:melt:Oberon0:core;
exports edu:umn:cs:melt:Oberon0:constructs:controlFlow;
exports edu:umn:cs:melt:Oberon0:constructs:procedures;

parser parse::Module_c {
  edu:umn:cs:melt:Oberon0:core;
  edu:umn:cs:melt:Oberon0:constructs:controlFlow;
  edu:umn:cs:melt:Oberon0:constructs:procedures;
}

