grammar edu:umn:cs:melt:Oberon0:tasks:lift:procedures;

imports edu:umn:cs:melt:Oberon0:core;
imports edu:umn:cs:melt:Oberon0:constructs:procedures;

imports edu:umn:cs:melt:Oberon0:tasks:lift:core;

imports silver:langutil;
imports silver:langutil:pp as pp;

