grammar edu:umn:cs:melt:Oberon0:core;

exports edu:umn:cs:melt:Oberon0:core:concreteSyntax;
exports edu:umn:cs:melt:Oberon0:core:abstractSyntax;

