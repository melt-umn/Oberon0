grammar edu:umn:cs:melt:Oberon0:components:L2;

exports edu:umn:cs:melt:Oberon0:core;
exports edu:umn:cs:melt:Oberon0:constructs:controlFlow;

parser parse::Module_c {
  edu:umn:cs:melt:Oberon0:core;
  edu:umn:cs:melt:Oberon0:constructs:controlFlow;
}


