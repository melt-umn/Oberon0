grammar edu:umn:cs:melt:exts:Oberon0:tables;

exports  edu:umn:cs:melt:exts:Oberon0:tables:concreteSyntax;