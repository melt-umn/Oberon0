grammar edu:umn:cs:melt:exts:silver:Oberon0;

exports edu:umn:cs:melt:exts:silver:Oberon0:concretesyntax;
