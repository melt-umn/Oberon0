grammar edu:umn:cs:melt:Oberon0:tasks:lift:dataStructures;

imports edu:umn:cs:melt:Oberon0:core;
imports edu:umn:cs:melt:Oberon0:constructs:dataStructures;

imports edu:umn:cs:melt:Oberon0:tasks:lift:core;


