grammar edu:umn:cs:melt:Oberon0:components:T3;

exports edu:umn:cs:melt:Oberon0:core:typeChecking;

