grammar edu:umn:cs:melt:Oberon0:components:L1;

exports edu:umn:cs:melt:Oberon0:core;

parser parse::Module_c {
  edu:umn:cs:melt:Oberon0:core;
}

