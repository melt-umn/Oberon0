grammar edu:umn:cs:melt:Oberon0:tasks:codegenC:procedures;

imports edu:umn:cs:melt:Oberon0:core;
imports edu:umn:cs:melt:Oberon0:constructs:procedures;

imports edu:umn:cs:melt:Oberon0:tasks:codegenC:core;

exports edu:umn:cs:melt:Oberon0:tasks:lift:procedures;

imports silver:langutil;
imports silver:langutil:pp as pp;

