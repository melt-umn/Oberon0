-- Control flow
grammar edu:umn:cs:melt:Oberon0:constructs:controlFlow;

{- exports both concrete and abstract syntax grammars to
   define the L2 extensions to L1. -}
exports edu:umn:cs:melt:Oberon0:constructs:controlFlow:concreteSyntax;
exports edu:umn:cs:melt:Oberon0:constructs:controlFlow:abstractSyntax;

