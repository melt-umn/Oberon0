grammar edu:umn:cs:melt:Oberon0:constructs:procedures;

exports edu:umn:cs:melt:Oberon0:constructs:procedures:abstractSyntax;
exports edu:umn:cs:melt:Oberon0:constructs:procedures:concreteSyntax;

